/*module Pong #(
	Y_SCREEN = 320,
	X_SCREEN = 240,
	MAX_SCORE = 10,
	BALL_SPEED,
	BALL_SIZE,
	PADDLE_SPEED,
	PADDLE_SIZE
	)(
	input clock,
	input reset,
	input start,
	input player1_up,
	input player1_down,
	input player2_up,
	input player2_down,
	);*/
//	
//	ClockDivider #(
//		CLOCK_IN		(50000000),
//		CLOCK_OUT	(4608000)
//		) PixelClock (
//		clk_in		(clock),
//		rst			(reset),
//		clk_out		()
//		)
		
	